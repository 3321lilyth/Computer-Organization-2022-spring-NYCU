`timescale 1ns/1ps
module MEMWB_register (
    input clk_i,
    input rst_i,
    input [3:0] WB_i,           //4 bit，MemToReg(拆成兩個WriteBack) 和 RegWite 和 jump
    input [31:0] DM_i,          //data memory 來的東西
    input [31:0] alu_ans_i,     //???????????????
    input [4:0] WBreg_i,        //rd    
    input [31:0] pc_add4_i,

    output reg [3:0] WB_o,
    output reg [31:0] DM_o,
    output reg [31:0] alu_ans_o,
    output reg [4:0] WBreg_o,
    output reg [31:0] pc_add4_o
);
/* Write your code HERE */
always @(posedge clk_i or negedge rst_i)begin
    if (~rst_i)begin //全部設定成0
        WB_o = 4'b0;
        DM_o = 32'b0;
        alu_ans_o = 32'b0;
        WBreg_o = 5'b0;
        pc_add4_o = 32'b0;
    end
    else begin
        WB_o = WB_i;
        DM_o = DM_i;
        alu_ans_o = alu_ans_i;
        WBreg_o = WBreg_i;
        pc_add4_o = pc_add4_i;
    end
    

end
endmodule
