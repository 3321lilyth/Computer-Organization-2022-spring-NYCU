`timescale 1ns/1ps
module Pipeline_CPU(
    clk_i,
    rst_i
);

//I/O port
input         clk_i;
input         rst_i;

//Internal Signals
wire [31:0] PC_i;
wire [31:0] PC_o;
wire [32-1:0] instr;
wire [31:0] MUXMemtoReg_o; //最後面要傳回來寫的資料之一
// wire [31:0] RD_data_Src;
wire [31:0] ALUResult;
// wire [31:0] MUXALUSrc_o;//?????有rs1、rs2，是哪一個拉幹
// wire [31:0] Decoder_o;
wire [31:0] RSdata_o;
wire [31:0] RTdata_o;
wire [31:0] Imm_Gen_o;
wire [32-1:0] Imm_4 = 4;
wire [31:0] ALUSrc1_3to1_o;
wire [31:0] ALUSrc2_3to1_o;
wire [31:0] ALUSrc2_2to1_o;
// wire [8:0]  MUX_control_o;

wire [31:0] PC_Add4;
wire [31:0] PC_Add_Immediate;

//控制
wire MUXControl;    // generated by hazard detection unit
wire PC_write;      // generated by hazard detection unit

wire [1:0] ALUOp;   // generated by main control
wire ALUSrc;
wire RegWrite;
wire Branch;
wire Jump;
wire WriteBackA, WriteBackB, MemRead, MemWrite;//MemtoReg 被我刪掉拆成兩個WriteBack了

wire Branch_zero;      //就是L2裡面的那個等號的 unit 吐出來的東西
wire PCSrc;
assign Branch_zero = (RSdata_o == RTdata_o )? 1:0;
assign PCSrc = Jump || (Branch && Branch_zero);

wire [31:0] ShiftLeft1_o; 
wire [31:0] DataMem_o;
wire [3:0] ALU_Ctrl_o;
wire ALU_zero;
wire [1:0] ForwardA;
wire [1:0] ForwardB;
wire [3:0] MUX_control_WB_o;
wire [1:0] MUX_control_Mem_o;
wire [2:0] MUX_control_Exe_o;

//Pipeline Register Signals
//IFID
wire [31:0] IFID_PC_o;
wire [31:0] IFID_Instr_o;
wire IFID_Write;
wire IFID_Flush;
assign IFID_Flush = Jump || (Branch && Branch_zero); //跟PCSrc 一模一樣
wire [31:0]IFID_PC_Add4_o;

//IDEXE
wire [31:0] IDEXE_Instr_o;
wire [3:0] IDEXE_WB_o;
wire [1:0] IDEXE_Mem_o;
wire [2:0] IDEXE_Exe_o;//L3，3 bit，{ALUOp,ALUSrc}
// wire [31:0] IDEXE_PC_o;
wire [31:0] IDEXE_RSdata_o;
wire [31:0] IDEXE_RTdata_o;
wire [31:0] IDEXE_ImmGen_o;
wire [3:0] IDEXE_Instr_30_14_12_o;
wire [31:0]IDEXE_PC_add4_o;
wire [4:0] IDEXE_RD_addr_o;
wire [4:0] IDEXE_RS1_addr_o;
wire [4:0] IDEXE_RS2_addr_o;

//EXEMEM
wire [31:0] EXEMEM_Instr_o; //不知為何要傳到L4的東西^^
wire [3:0] EXEMEM_WB_o;
wire [1:0] EXEMEM_Mem_o;//2 bit，{MemRead,MemWrite}，沒有 branch因為 branch 移到L2了
// wire [31:0] EXEMEM_PCsum_o;
wire EXEMEM_Zero_o;//不知為何要傳到L4的東西^^
wire [31:0] EXEMEM_ALUResult_o;
wire [31:0] EXEMEM_RTdata_o;
wire [4:0]  EXEMEM_RD_addr_o;
wire [31:0] EXEMEM_PC_Add4_o;

//MEMWB
wire [3:0] MEMWB_WB_o; //4 bit，{RegWrite,WriteBackA,WriteBackB,jump}
wire [31:0] MEMWB_DM_o;
wire [31:0] MEMWB_ALUresult_o;
wire [4:0]  MEMWB_RD_addr_o;
wire [31:0] MEMWB_PC_Add4_o;//不知為何要傳到L5的東西^^

wire debug;

assign debug = 0;

// IF
MUX_2to1 MUX_PCSrc(
    .data0_i(PC_Add4),
    .data1_i(PC_Add_Immediate),
    .select_i(PCSrc),
    .data_o(PC_i)
    
);

ProgramCounter PC(
    .clk_i(clk_i),
    .rst_i(rst_i),
    .PCWrite(PC_write),//PC_write
    .pc_i(PC_i),
    .pc_o(PC_o)
);

Adder PC_plus_4_Adder(
    .src1_i(PC_o),
    .src2_i(Imm_4),
    .sum_o(PC_Add4)

);

Instr_Memory IM(
    .addr_i(PC_o), //32
    .instr_o(instr) //32
);

IFID_register IFtoID(
    .clk_i(clk_i),
    .rst_i(rst_i),
    .flush(IFID_Flush),
    .IFID_write(IFID_Write),
    .address_i(PC_o),
    .instr_i(instr),
    .pc_add4_i(PC_Add4),

    .address_o(IFID_PC_o),
    .instr_o(IFID_Instr_o),
    .pc_add4_o(IFID_PC_Add4_o)
);

// ID

Hazard_detection Hazard_detection_obj(
    .IFID_regRs(IFID_Instr_o[19:15]),
    .IFID_regRt(IFID_Instr_o[24:20]),
    .IDEXE_regRd(IDEXE_RD_addr_o),
    .IDEXE_memRead(IDEXE_Mem_o[1]),

    .PC_write(PC_write),
    .IFID_write(IFID_Write),
    .control_output_select(MUXControl) 
);
// assign WB_i[0] = Jump;
// assign WB_i[1] = WriteBackB;
// assign WB_i[2] = WriteBackA;
// assign WB_i[3] = RegWrite;

wire [1:0] tmp;
assign tmp = {MemRead,MemWrite};
wire [3:0] WB_i;
assign WB_i = {RegWrite,WriteBackA,WriteBackB,Jump};
MUX_control MUX_control( //ID/EX 三個 control 前面的那個 MUX
    .WB_i(WB_i),        //4 bit，RegWite 和 MemToReg(拆成{WriteBackA}{WriteBackB}) {jump}
    .Mem_i({MemRead,MemWrite}),       //2 bit，{MemRead}{MemWrite}，沒有 branch因為 branch 移到L2了
    .Exe_i({ALUOp,ALUSrc}),       //L3，3 bit，{ALU op*2}{ALU_src}
    .hazard_control(MUXControl),

    //output
    .WB_o(MUX_control_WB_o),
    .Mem_o(MUX_control_Mem_o),
    .Exe_o(MUX_control_Exe_o)

);

Decoder Decoder(
    .instr_i(IFID_Instr_o),

    .RegWrite(RegWrite),
    .Branch(Branch),
    .Jump(Jump),
    .MemRead(MemRead),
    .MemWrite(MemWrite),

    .WriteBackA(WriteBackA),    
    .WriteBackB(WriteBackB),
    .ALUSrc(ALUSrc),
    .ALUOp(ALUOp)
);

// MUX_2to1 MUX_RD_data_Src(//有沒有可能先用了上次的 jump 然後這次的 decoder 才解出這次的 jump
//     .data0_i(MUXMemtoReg_o),
//     .data1_i(IFID_PC_Add4_o),
//     .select_i(Jump),
//     .data_o(RD_data_Src)
// );

Reg_File RF(
    .clk_i(clk_i),
    .rst_i(rst_i),
    .RSaddr_i(IFID_Instr_o[19:15]),
    .RTaddr_i(IFID_Instr_o[24:20]),
    .RDaddr_i(MEMWB_RD_addr_o),
    .RDdata_i(MUXMemtoReg_o),

    .RegWrite_i(MEMWB_WB_o[3]), //MEMWB_WB_o[3]

    .RSdata_o(RSdata_o),
    .RTdata_o(RTdata_o)
);

Imm_Gen ImmGen(
    .instr_i(IFID_Instr_o),
    .Imm_Gen_o(Imm_Gen_o)
);

Shift_Left_1 SL1(
    .data_i(Imm_Gen_o),
    .data_o(ShiftLeft1_o)
);

Adder Branch_Adder(
    .src1_i(IFID_PC_o),
    .src2_i(ShiftLeft1_o),
    .sum_o(PC_Add_Immediate)
);

IDEXE_register IDtoEXE(
    .clk_i(clk_i),
    .rst_i(rst_i),
    .instr_i(IFID_Instr_o),
    
    .WB_i(MUX_control_WB_o),
    .Mem_i(MUX_control_Mem_o),
    .Exe_i(MUX_control_Exe_o),
    .data1_i(RSdata_o),
    .data2_i(RTdata_o),

    .immgen_i(Imm_Gen_o),
    .alu_ctrl_instr({IFID_Instr_o[30],IFID_Instr_o[14:12]}),
    .WBreg_i(IFID_Instr_o[11:7]),
    .pc_add4_i(IFID_PC_Add4_o),
    .RS1_i(IFID_Instr_o[19:15]),
    .RS2_i(IFID_Instr_o[24:20]),
    
    //output
    .instr_o(IDEXE_Instr_o),
    .WB_o(IDEXE_WB_o),
    .Mem_o(IDEXE_Mem_o),
    .Exe_o(IDEXE_Exe_o),
    
    .data1_o(IDEXE_RSdata_o),
    .data2_o(IDEXE_RTdata_o),
    .immgen_o(IDEXE_ImmGen_o),
    .alu_ctrl_input(IDEXE_Instr_30_14_12_o),
    .WBreg_o(IDEXE_RD_addr_o),
    .pc_add4_o(IDEXE_PC_add4_o),
    .RS1_o(IDEXE_RS1_addr_o),
    .RS2_o(IDEXE_RS2_addr_o)
);

// EXE
MUX_2to1 MUX_ALUSrc(
    .data0_i(ALUSrc2_3to1_o),
    .data1_i(IDEXE_ImmGen_o),
    .select_i(IDEXE_Exe_o[0]),
    .data_o(ALUSrc2_2to1_o)
);

ForwardingUnit FWUnit(
    .IDEXE_RS1(IDEXE_RS1_addr_o),
    .IDEXE_RS2(IDEXE_RS2_addr_o),
    .EXEMEM_RD(EXEMEM_RD_addr_o),
    .MEMWB_RD(MEMWB_RD_addr_o),
    .EXEMEM_RegWrite(EXEMEM_WB_o[3]),
    .MEMWB_RegWrite(MEMWB_WB_o[3]),

    //output
    .ForwardA(ForwardA),
    .ForwardB(ForwardB)
);

MUX_3to1 MUX_ALU_src1(
    .data0_i(IDEXE_RSdata_o),
    .data1_i(MUXMemtoReg_o),
    .data2_i(EXEMEM_ALUResult_o),
    .select_i(ForwardA),
    .data_o(ALUSrc1_3to1_o)
);

MUX_3to1 MUX_ALU_src2(
    .data0_i(IDEXE_RTdata_o),
    .data1_i(MUXMemtoReg_o),
    .data2_i(EXEMEM_ALUResult_o),
    .select_i(ForwardB),
    .data_o(ALUSrc2_3to1_o)
);

ALU_Ctrl ALU_Ctrl(
    .instr(IDEXE_Instr_30_14_12_o),
    .ALUOp(IDEXE_Exe_o[2:1]),
    .ALU_Ctrl_o(ALU_Ctrl_o)
);

alu alu(
    .rst_n(rst_i),
    .src1(ALUSrc1_3to1_o),
    .src2(ALUSrc2_2to1_o),
    .ALU_control(ALU_Ctrl_o),
    .result(ALUResult),
    .zero(ALU_zero)
);

EXEMEM_register EXEtoMEM(
    .clk_i(clk_i),
    .rst_i(rst_i),
    .instr_i(IDEXE_Instr_o),
    .WB_i(IDEXE_WB_o),
    .Mem_i(IDEXE_Mem_o),
    .zero_i(ALU_zero),
    .alu_ans_i(ALUResult),
    .rtdata_i(ALUSrc2_3to1_o),
    .WBreg_i(IDEXE_RD_addr_o),
    .pc_add4_i(IDEXE_PC_add4_o),
    
    //output
    .instr_o(EXEMEM_Instr_o),
    .WB_o(EXEMEM_WB_o),
    .Mem_o(EXEMEM_Mem_o),
    .zero_o(EXEMEM_Zero_o),
    .alu_ans_o(EXEMEM_ALUResult_o),
    .rtdata_o(EXEMEM_RTdata_o),
    .WBreg_o(EXEMEM_RD_addr_o),
    .pc_add4_o(EXEMEM_PC_Add4_o)
);

// MEM
Data_Memory Data_Memory(
    .clk_i(clk_i),
    .addr_i(EXEMEM_ALUResult_o),
    .data_i(EXEMEM_RTdata_o),
    .MemRead_i(EXEMEM_Mem_o[1]),
    .MemWrite_i(EXEMEM_Mem_o[0]),
    .data_o(DataMem_o)
);

MEMWB_register MEMtoWB(
    .clk_i(clk_i),
    .rst_i(rst_i),
    .WB_i(EXEMEM_WB_o),
    .DM_i(DataMem_o),
    .alu_ans_i(EXEMEM_ALUResult_o),
    .WBreg_i(EXEMEM_RD_addr_o),
    .pc_add4_i(EXEMEM_PC_Add4_o),

    //output
    .WB_o(MEMWB_WB_o),
    .DM_o(MEMWB_DM_o),
    .alu_ans_o(MEMWB_ALUresult_o),
    .WBreg_o(MEMWB_RD_addr_o),
    .pc_add4_o(MEMWB_PC_Add4_o)
);

wire [31:0] MUX_MemtoReg_o;
// WB
MUX_2to1 MUX_MemtoReg(
    .data0_i(MEMWB_DM_o),
    .data1_i(MEMWB_ALUresult_o),
    .select_i(MEMWB_WB_o[2]),
    .data_o(MUX_MemtoReg_o)

);

MUX_2to1 MUX_jump(
    .data0_i(MUX_MemtoReg_o),
    .data1_i(MEMWB_PC_Add4_o),
    .select_i(MEMWB_WB_o[0]),
    .data_o(MUXMemtoReg_o)

);

endmodule



